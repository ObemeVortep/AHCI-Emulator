/*
 * Global debug configuration flags:
 * 
 * - Enables USB-based debug output path and conditionally activates internal diagnostic modules.
 * - Each define toggles logging and inspection for a specific subsystem or dataflow.
 * - Designed for modular debugging with strict dependency on a central debug interface flag.
 * - Requires corresponding Vivado IP blocks to be manually disabled when the main flag is inactive.
 * 
 * Code has been redacted for ethical and security reasons.
 * 22 LOC
 */
/*
 * Module responsible for providing SMART data sectors of the disk.
 *
 * Stores the device's SMART data structure in block RAM and delivers it on read requests.
 *
 * Code has been redacted for ethical and security reasons.
 * 44 LOC
 */
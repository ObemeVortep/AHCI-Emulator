/*
 * This module coordinates the monitoring process by managing data flow and control signals:
 *
 * - Operates after required initializations and address resolutions.
 * - Receives base addresses needed for data access.
 * - Controls two submodules: a main controller handling data parsing and a helper managing PCIe transactions.
 * - Handles virtual address reads and data retrieval through these submodules.
 * - Continuously processes and outputs updated data once initialized.
 *
 * Code has been redacted for ethical and security reasons.
 * 143 LOC
 */
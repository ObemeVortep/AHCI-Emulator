/*
 * Configuration header defining scanning granularity and memory bounds:
 * 
 * - Selects memory read length for scan operations via mutually exclusive macros.
 * - Sets associated constants for each scan mode:
 *     - Read request length.
 *     - Byte enable mask.
 *     - Address increment and alignment constraints.
 *     - Bit width reduction for analyzer logic.
 * - Specifies total physical memory size to bound scanning region.
 * - Provides consistent constants for scanner and analyzer modules.
 * 
 * Code has been redacted for ethical and security reasons.
 * 83 LOC
 */